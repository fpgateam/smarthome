  --Example instantiation for system 'lcd'
  lcd_inst : lcd
    port map(
      LCD_E_from_the_lcd_0 => LCD_E_from_the_lcd_0,
      LCD_RS_from_the_lcd_0 => LCD_RS_from_the_lcd_0,
      LCD_RW_from_the_lcd_0 => LCD_RW_from_the_lcd_0,
      LCD_data_to_and_from_the_lcd_0 => LCD_data_to_and_from_the_lcd_0,
      out_port_from_the_pio_0 => out_port_from_the_pio_0,
      clk_0 => clk_0,
      reset_n => reset_n
    );


